// alu option
`define ALU_OP_WD   11
`define ALU_ADD     0
`define ALU_SUB     1
`define ALU_SLT     2
`define ALU_SLTU    3
`define ALU_XOR     4
`define ALU_OR      5
`define ALU_AND     6
`define ALU_SLL     7
`define ALU_SRL     8
`define ALU_SRA     9
`define ALU_LUI     10
// bus size
`define F_TO_D_BUS_WD  64
`define D_TO_E_BUS_WD  163
`define E_TO_M_BUS_WD  107
`define M_TO_W_BUS_WD  103
`define W_TO_RF_BUS_WD 38
`define D_TO_H_BUS_WD  12
`define E_TO_H_BUS_WD  17
`define M_TO_H_BUS_WD  7
`define W_TO_H_BUS_WD  6